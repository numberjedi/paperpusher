version https://git-lfs.github.com/spec/v1
oid sha256:3aff8bd2ea50bc4cb88b8a1b64071929a20a49a72dccf5200e7aa54a9e3ee992
size 712
